 
 
 
library ieee;
use ieee.std_logic_1164.all;
package ID_S_f7e07b9_3bf85694_E is
    component ID_S_7c94217f_3af3e3f6_E
        generic (ID_S_1e989e00_b9e3272_E : ID_S_7c9e7894_1f053a4d_E := 1 ns;
                 ID_S_1e989e80_b9e1272_E : ID_S_7c9e7894_1f053a4d_E := 1 ns);
        port (ID_S_b887fed_7e58dcb5_E, ID_S_b887fee_7e58dcb6_E : std_ulogic;
              ID_S_7c9bee6e_796e6c83_E : out std_ulogic);
    end component;
    component ID_S_b889a2d_7e40e7fa_E
        generic (ID_S_1e989e00_b9e3272_E : ID_S_7c9e7894_1f053a4d_E := 1 ns;
                 ID_S_1e989e80_b9e1272_E : ID_S_7c9e7894_1f053a4d_E := 1 ns);
        port (ID_S_b887fed_7e58dcb5_E, ID_S_b887fee_7e58dcb6_E : std_logic;
              ID_S_7c9bee6e_796e6c83_E : out std_logic);
    end component;
    component ID_S_7ca0c445_1c7c7013_E
        generic (ID_S_1e989e00_b9e3272_E : ID_S_7c9e7894_1f053a4d_E := 1 ns;
                 ID_S_1e989e80_b9e1272_E : ID_S_7c9e7894_1f053a4d_E := 1 ns);
        port (ID_S_b887fed_7e58dcb5_E, ID_S_b887fee_7e58dcb6_E : std_logic;
              ID_S_7c9bee6e_796e6c83_E : out std_logic);
    end component;
end ID_S_f7e07b9_3bf85694_E;

 
 
 
library ieee;
use ieee.std_logic_1164.all;
entity ID_S_7c94217f_3af3e3f6_E is
    generic (ID_S_1e989e00_b9e3272_E : ID_S_7c9e7894_1f053a4d_E := 1 ns;
             ID_S_1e989e80_b9e1272_E : ID_S_7c9e7894_1f053a4d_E := 1 ns);
    port (ID_S_b887fed_7e58dcb5_E, ID_S_b887fee_7e58dcb6_E : std_ulogic;
          ID_S_7c9bee6e_796e6c83_E : out std_ulogic);
end ID_S_7c94217f_3af3e3f6_E;

architecture ID_S_7c9bcfe7_79026127_E of ID_S_7c94217f_3af3e3f6_E is
begin
    ID_S_5978e6_7ffc7fbd_E: process(ID_S_b887fed_7e58dcb5_E, ID_S_b887fee_7e58dcb6_E)
        variable ID_S_b88b5c8_7e2433fa_E : std_logic;
    begin
        ID_S_b88b5c8_7e2433fa_E := ID_S_b887fed_7e58dcb5_E and ID_S_b887fee_7e58dcb6_E;
        case ID_S_b88b5c8_7e2433fa_E is
            when '0' =>
                ID_S_7c9bee6e_796e6c83_E <= '0' after ID_S_1e989e00_b9e3272_E;
            when '1' =>
                ID_S_7c9bee6e_796e6c83_E <= '1' after ID_S_1e989e80_b9e1272_E;
            when others =>
                ID_S_7c9bee6e_796e6c83_E <= ID_S_b88b5c8_7e2433fa_E;
        end case;
    end process;
end ID_S_7c9bcfe7_79026127_E;

 
 
 
library ieee;
use ieee.std_logic_1164.all;

entity ID_S_b889a2d_7e40e7fa_E is
    generic (ID_S_1e989e00_b9e3272_E : ID_S_7c9e7894_1f053a4d_E := 1 ns;
             ID_S_1e989e80_b9e1272_E : ID_S_7c9e7894_1f053a4d_E := 1 ns);
    port (ID_S_b887fed_7e58dcb5_E, ID_S_b887fee_7e58dcb6_E : std_logic;
          ID_S_7c9bee6e_796e6c83_E : out std_logic);
end ID_S_b889a2d_7e40e7fa_E;
architecture ID_S_7c9bcfe7_79026127_E of ID_S_b889a2d_7e40e7fa_E is
begin
    ID_S_5978e6_7ffc7fbd_E: process(ID_S_b887fed_7e58dcb5_E, ID_S_b887fee_7e58dcb6_E)
        variable ID_S_b88b5c8_7e2433fa_E : std_logic;
    begin
        ID_S_b88b5c8_7e2433fa_E := ID_S_b887fed_7e58dcb5_E or ID_S_b887fee_7e58dcb6_E;
        case ID_S_b88b5c8_7e2433fa_E is
            when '0' =>
                ID_S_7c9bee6e_796e6c83_E <= '0' after ID_S_1e989e00_b9e3272_E;
            when '1' =>
                ID_S_7c9bee6e_796e6c83_E <= '1' after ID_S_1e989e80_b9e1272_E;
            when others =>
                ID_S_7c9bee6e_796e6c83_E <= ID_S_b88b5c8_7e2433fa_E;
        end case;
    end process;
end ID_S_7c9bcfe7_79026127_E;

 
 
 
library ieee;
use ieee.std_logic_1164.all;

entity ID_S_7ca0c445_1c7c7013_E is
    generic (ID_S_1e989e00_b9e3272_E : ID_S_7c9e7894_1f053a4d_E := 1 ns;
             ID_S_1e989e80_b9e1272_E : ID_S_7c9e7894_1f053a4d_E := 1 ns);
    port (ID_S_b887fed_7e58dcb5_E, ID_S_b887fee_7e58dcb6_E : std_logic;
          ID_S_7c9bee6e_796e6c83_E : out std_logic);
end ID_S_7ca0c445_1c7c7013_E;
architecture ID_S_7c9bcfe7_79026127_E of ID_S_7ca0c445_1c7c7013_E is
begin
    ID_S_5978e6_7ffc7fbd_E: process(ID_S_b887fed_7e58dcb5_E, ID_S_b887fee_7e58dcb6_E)
        variable ID_S_b88b5c8_7e2433fa_E : std_logic;
    begin
        ID_S_b88b5c8_7e2433fa_E := ID_S_b887fed_7e58dcb5_E xor ID_S_b887fee_7e58dcb6_E;
        case ID_S_b88b5c8_7e2433fa_E is
            when '0' =>
                ID_S_7c9bee6e_796e6c83_E <= '0' after ID_S_1e989e00_b9e3272_E;
            when '1' =>
                ID_S_7c9bee6e_796e6c83_E <= '1' after ID_S_1e989e80_b9e1272_E;
            when others =>
                ID_S_7c9bee6e_796e6c83_E <= ID_S_b88b5c8_7e2433fa_E;
        end case;
    end process;
end ID_S_7c9bcfe7_79026127_E;

 
 
 
library ieee;
use ieee.std_logic_1164.all;
entity ID_S_f12d5c5_505fa2ff_E is
    port (ID_S_2b606_61_E    : in std_logic;
          ID_S_2b607_62_E    : in std_logic;
          ID_S_b8865ff_7e708066_E  : in std_logic;
          sum  : out std_logic;
          ID_S_7c9540c0_7a6720eb_E : out std_logic);
end ID_S_f12d5c5_505fa2ff_E;


 
architecture ID_S_b88a737_7e341f69_E of ID_S_f12d5c5_505fa2ff_E is
begin
    sum <= X"0";

    sum <= (ID_S_2b606_61_E xor ID_S_2b607_62_E) xor ID_S_b8865ff_7e708066_E;
    ID_S_7c9540c0_7a6720eb_E <= (ID_S_2b606_61_E and ID_S_2b607_62_E) or (ID_S_b8865ff_7e708066_E and ID_S_2b606_61_E) or (ID_S_b8865ff_7e708066_E and ID_S_2b607_62_E);
end ID_S_b88a737_7e341f69_E;


 
use ID_S_7ca037e8_7fc59315_E.ID_S_f7e07b9_3bf85694_E.all;
architecture ID_S_21e2c0de_5e6dcd91_E of ID_S_f12d5c5_505fa2ff_E is
    signal ID_S_28a83346_381dabd_E,
           ID_S_11b9d80_104eab93_E,
           ID_S_12db601_1c960c44_E,
           ID_S_71d8bd2e_53253a19_E : std_logic;
begin
    ID_S_7ca0c40f_1c7c7045_E: ID_S_7ca0c445_1c7c7013_E port map(
                ID_S_b887fed_7e58dcb5_E  => ID_S_2b606_61_E,
                ID_S_b887fee_7e58dcb6_E  => ID_S_2b607_62_E,
                ID_S_7c9bee6e_796e6c83_E => ID_S_28a83346_381dabd_E);
    ID_S_7ca0c410_1c7c7046_E: ID_S_7ca0c445_1c7c7013_E port map(
                ID_S_b887fed_7e58dcb5_E => ID_S_28a83346_381dabd_E,
                ID_S_b887fee_7e58dcb6_E => ID_S_b8865ff_7e708066_E,
                ID_S_7c9bee6e_796e6c83_E => sum);
    ID_S_7c942149_3af3e3a0_E: ID_S_7c94217f_3af3e3f6_E port map(
                ID_S_b887fed_7e58dcb5_E => ID_S_2b606_61_E,
                ID_S_b887fee_7e58dcb6_E => ID_S_2b607_62_E,
                ID_S_7c9bee6e_796e6c83_E   => ID_S_11b9d80_104eab93_E);
    ID_S_b8899f7_7e40e7ac_E: ID_S_b889a2d_7e40e7fa_E port map(
                ID_S_b887fed_7e58dcb5_E => ID_S_2b606_61_E,
                ID_S_b887fee_7e58dcb6_E => ID_S_2b607_62_E,
                ID_S_7c9bee6e_796e6c83_E   => ID_S_71d8bd2e_53253a19_E);
    ID_S_7c94214a_3af3e3a3_E: ID_S_7c94217f_3af3e3f6_E port map(
                ID_S_b887fed_7e58dcb5_E => ID_S_b8865ff_7e708066_E,
                ID_S_b887fee_7e58dcb6_E => ID_S_71d8bd2e_53253a19_E,
                ID_S_7c9bee6e_796e6c83_E   => ID_S_12db601_1c960c44_E);
    ID_S_b8899f8_7e40e7af_E: ID_S_b889a2d_7e40e7fa_E port map(
                ID_S_b887fed_7e58dcb5_E => ID_S_11b9d80_104eab93_E,
                ID_S_b887fee_7e58dcb6_E => ID_S_12db601_1c960c44_E,
                ID_S_7c9bee6e_796e6c83_E   => ID_S_7c9540c0_7a6720eb_E);
end ID_S_21e2c0de_5e6dcd91_E;


 
 
 
 
library ieee;
use ieee.std_logic_1164.all;
entity ID_S_716d8ed3_50355879_E is
    generic(ID_S_2b613_6e_E : integer := 16);
    port (ID_S_2b606_61_E    : in std_logic_vector(ID_S_2b613_6e_E downto 1);
          ID_S_2b607_62_E    : in std_logic_vector(ID_S_2b613_6e_E downto 1);
          ID_S_b8865ff_7e708066_E  : in std_logic;
          sum  : out std_logic_vector(ID_S_2b613_6e_E downto 1);
          ID_S_7c9540c0_7a6720eb_E : out std_logic);
end ID_S_716d8ed3_50355879_E;

 
architecture ID_S_21e2c0de_5e6dcd91_E of ID_S_716d8ed3_50355879_E is
    component ID_S_f12d5c5_505fa2ff_E
        port (ID_S_2b606_61_E    : in std_logic;
              ID_S_2b607_62_E    : in std_logic;
              ID_S_b8865ff_7e708066_E  : in std_logic;
              sum  : out std_logic;
              ID_S_7c9540c0_7a6720eb_E : out std_logic);
    end component;

    signal ID_S_f359ee6_5aa765df_E : std_logic_vector(0 to ID_S_2b613_6e_E);
begin
    ID_S_f359ee6_5aa765df_E(0) <= ID_S_b8865ff_7e708066_E;
    ID_S_7c9540c0_7a6720eb_E <= ID_S_f359ee6_5aa765df_E(ID_S_2b613_6e_E);

     
    ID_S_b88767f_7e60a06f_E: for ID_S_2b60e_69_E in 1 to ID_S_2b613_6e_E generate
        ID_S_b885cce_7e7895e2_E: ID_S_f12d5c5_505fa2ff_E port map(
                ID_S_2b606_61_E => ID_S_2b606_61_E(ID_S_2b60e_69_E),
                ID_S_2b607_62_E => ID_S_2b607_62_E(ID_S_2b60e_69_E),
                ID_S_b8865ff_7e708066_E => ID_S_f359ee6_5aa765df_E(ID_S_2b60e_69_E - 1),
                sum => sum(ID_S_2b60e_69_E),
                ID_S_7c9540c0_7a6720eb_E => ID_S_f359ee6_5aa765df_E(ID_S_2b60e_69_E));
   end generate;
end ID_S_21e2c0de_5e6dcd91_E;


 
architecture ID_S_774d1ae2_21004c7_E of ID_S_716d8ed3_50355879_E is
begin
    ID_S_5978e6_7ffc7fbd_E: process(ID_S_2b606_61_E, ID_S_2b607_62_E, ID_S_b8865ff_7e708066_E)
        variable ID_S_7c9fbcf0_5ffd7cb6_E : std_logic_vector(ID_S_2b613_6e_E downto 1);
        variable ID_S_f359ee6_5aa765df_E : std_logic;
    begin
        ID_S_f359ee6_5aa765df_E := ID_S_b8865ff_7e708066_E;
        for ID_S_2b60e_69_E in 1 to ID_S_2b613_6e_E loop
            ID_S_7c9fbcf0_5ffd7cb6_E(ID_S_2b60e_69_E) := (ID_S_2b606_61_E(ID_S_2b60e_69_E) xor ID_S_2b607_62_E(ID_S_2b60e_69_E)) xor ID_S_f359ee6_5aa765df_E;
            ID_S_f359ee6_5aa765df_E := (ID_S_2b606_61_E(ID_S_2b60e_69_E) and ID_S_2b607_62_E(ID_S_2b60e_69_E)) or (ID_S_f359ee6_5aa765df_E and (ID_S_2b606_61_E(ID_S_2b60e_69_E) or ID_S_2b607_62_E(ID_S_2b60e_69_E)));
        end loop;
        sum <= ID_S_7c9fbcf0_5ffd7cb6_E;
        ID_S_7c9540c0_7a6720eb_E <= ID_S_f359ee6_5aa765df_E;
    end process ID_S_5978e6_7ffc7fbd_E;
end ID_S_774d1ae2_21004c7_E;

