   module ID_S_56f8898b_39580807_E  (    input1,  ID_S_597800_7ffcb7a7_E,    ID_S_5978c5_7ffc87a2_E,  ID_S_5978c6_7ffc87a1_E  );      input input1;  input ID_S_597800_7ffcb7a7_E;      output ID_S_5978c5_7ffc87a2_E;  output ID_S_5978c6_7ffc87a1_E;    assign ID_S_5978c5_7ffc87a2_E = input1 & ID_S_597800_7ffcb7a7_E;  assign ID_S_5978c6_7ffc87a1_E = ^{input1,ID_S_597800_7ffcb7a7_E};    endmodule   